ENTITY MARCAPASSO IS
  PORT(
  RESET,SENSORA,SENSORV,CLK_IN:IN BIT;
  TEMPOA: IN INTEGER RANGE 0 TO 15;
  TEMPOV: IN INTEGER RANGE 0 TO 15;
  OUT_PA,OUT_PV: OUT BIT;
  SAIDA_DISPA:OUT BIT_VECTOR(6 DOWNTO 0);--A..G
  ENABLE_DISPA,ENABLE_DISPV:OUT BIT);
END MARCAPASSO;

ARCHITECTURE ONE OF MARCAPASSO IS
  COMPONENT MAQESTADO
    PORT(
    CLK,RESET,SENSORA,SENSORV,TIMEA,TIMEV: IN BIT;
    ENABLEA,ENABLEV,OUT_PA,OUT_PV: OUT BIT);
  END COMPONENT;

  COMPONENT DIV_CLK
    PORT(
    RESET,CLK_IN: IN BIT;
    CLK_OUT1: OUT BIT;
    CLK_OUT2: OUT BIT);
  END COMPONENT;

  COMPONENT TIMER
    PORT(
    CLK,ENABLE,RESET: IN BIT;
    TEMPO: IN INTEGER RANGE 0 TO 15;
    SAIDA: OUT BIT);
  END COMPONENT;

  COMPONENT CONT_DEC
    PORT(
    IN_CONT,RESET: IN BIT;
    SAIDA_DISP: OUT BIT_VECTOR(6 DOWNTO 0));--A..G
  END COMPONENT;

  COMPONENT MUX
    PORT(
          CLK: IN BIT;
    DISPA,DISPV: IN BIT_VECTOR(6 DOWNTO 0);
    SAIDA_DISP: OUT BIT_VECTOR(6 DOWNTO 0);--A..G
    ENABLE_DISPA,ENABLE_DISPV:OUT BIT);
  END COMPONENT;

  SIGNAL X1,X2,X3,X4,X5,X6,X7,X8,X9,X10:BIT;
  SIGNAL Y1,Y2:BIT_VECTOR(6 DOWNTO 0);
BEGIN
  CHIP1: DIV_CLK PORT MAP (RESET=>RESET,CLK_IN=>CLK_IN,CLK_OUT1=>X1,CLK_OUT2=>X10);
  CHIP2: MAQESTADO PORT MAP (CLK=>X1,RESET=>RESET,SENSORA=>SENSORA,SENSORV=>SENSORV,
                             TIMEA=>X2,TIMEV=>X3,ENABLEA=>X4,ENABLEV=>X5,OUT_PA=>X8,OUT_PV=>X9);
  CHIP3: TIMER PORT MAP (CLK=>X1,ENABLE=>X5,TEMPO=>TEMPOV,SAIDA=>X3,RESET=>RESET);
  CHIP4: TIMER PORT MAP (CLK=>X1,ENABLE=>X4,TEMPO=>TEMPOA,SAIDA=>X2,RESET=>RESET);
  CHIP5: CONT_DEC PORT MAP (IN_CONT=>X8,RESET=>RESET,SAIDA_DISP=>Y1);
  CHIP6: CONT_DEC PORT MAP (IN_CONT=>X9,RESET=>RESET,SAIDA_DISP=>Y2);
  CHIP7: MUX PORT MAP (CLK=>X10,DISPA=>Y1,DISPV=>Y2,SAIDA_DISP=>SAIDA_DISPA,ENABLE_DISPA=>ENABLE_DISPA,
                       ENABLE_DISPV=>ENABLE_DISPV);
  OUT_PA<=X8;
  OUT_PV<=X9;
END ONE;

ENTITY MAQESTADO IS
  PORT(
  CLK,RESET,SENSORA,SENSORV,TIMEA,TIMEV: IN BIT;
  ENABLEA,ENABLEV,OUT_PA,OUT_PV: OUT BIT);
END MAQESTADO;

ARCHITECTURE ONE OF MAQESTADO IS
  TYPE STATE IS (WAITV,WAITA,PA,PV);
  SIGNAL X: STATE;
BEGIN
  PROCESS (CLK)
  BEGIN 
    IF RESET='0'THEN
      X<=WAITV;

    ELSIF CLK'EVENT AND CLK='1'THEN
      CASE X IS
        WHEN WAITV => --X<=PV;
          IF TIMEV='1' THEN X<=PV;
          ELSIF SENSORV='0'THEN X<= WAITA;
          END IF;
        WHEN WAITA =>-- X<=PA;
          IF TIMEA='1' THEN X<=PA;
          ELSIF SENSORA='0'THEN X<= WAITV;
          END IF;
        WHEN PA =>
          X<= WAITV;
        WHEN PV =>
          X<= WAITA;
      END CASE;
    END IF;
  END PROCESS;
  WITH X SELECT
    OUT_PA<='1' WHEN PA,
            '0' WHEN PV,
            '0' WHEN WAITA,
            '0' WHEN WAITV;

  WITH X SELECT
    OUT_PV <='1' WHEN PV,
             '0' WHEN PA,
             '0' WHEN WAITA,
             '0' WHEN WAITV;	
  WITH X SELECT
    ENABLEA <='0' WHEN PV,
              '0' WHEN PA,
              '1' WHEN WAITA,
              '0' WHEN WAITV;			  
  WITH X SELECT
    ENABLEV <='0' WHEN PV,
              '0' WHEN PA,
              '0' WHEN WAITA,
              '1' WHEN WAITV;   


END ONE;

ENTITY DIV_CLK IS
  PORT(
  RESET,CLK_IN: IN BIT;
  CLK_OUT1: OUT BIT;
  CLK_OUT2: OUT BIT);
END DIV_CLK;

ARCHITECTURE ONE OF DIV_CLK IS
  SIGNAL X:INTEGER RANGE 0 TO 2500000;
  SIGNAL X1:INTEGER RANGE 0 TO 2500000;

  SIGNAL AUX:BIT:='0';
  SIGNAL AUX1:BIT:='0';

BEGIN
  PROCESS (CLK_IN,reset)
  BEGIN 
    IF RESET='0'THEN
      X<=0;
      X1<=0;		
    ELSIF CLK_IN'EVENT AND CLK_IN='1'THEN
      IF X=2500000  THEN 
        X<=0;
        AUX<=NOT AUX;
      ELSE
        X<=X+1;
      END IF;
      IF X1=25000  THEN 
        X1<=0;
        AUX1<=NOT AUX1;
      ELSE
        X1<=X1+1;
      END IF;
    END IF;
  END PROCESS;
  CLK_OUT1<=AUX;
  CLK_OUT2<=AUX1;
END ONE;

ENTITY TIMER IS
  PORT(
  CLK,ENABLE,RESET: IN BIT;
  TEMPO: IN INTEGER RANGE 0 TO 15;
  SAIDA: OUT BIT);
END TIMER;
ARCHITECTURE ONE OF TIMER IS
  SIGNAL X: INTEGER RANGE 0 TO 15;
BEGIN
  PROCESS (CLK,RESET)
  BEGIN 
    IF  RESET='0'THEN
      X<=TEMPO;
      SAIDA<='0';
    ELSIF CLK'EVENT AND CLK='1'THEN
      IF ENABLE='0'THEN
        X<=TEMPO;
        SAIDA<='0'; 
      ELSIF (X=0) AND (ENABLE='1') THEN 
        SAIDA<='1';
      ELSIF (X>0) AND (ENABLE='1') THEN
        X<=X-1;
        SAIDA<='0'; 
      END IF;
    END IF;
  END PROCESS;
END ONE;
ENTITY CONT_DEC IS
  PORT(
  IN_CONT,RESET: IN BIT;
  SAIDA_DISP: OUT BIT_VECTOR(6 DOWNTO 0));--A..G
END CONT_DEC;

ARCHITECTURE ONE OF CONT_DEC IS
  SIGNAL X: INTEGER RANGE 0 TO 9;
BEGIN
  PROCESS (IN_CONT,RESET)
  BEGIN 
    IF  RESET='0'THEN
      X<= 0;
    ELSIF IN_CONT'EVENT AND IN_CONT='1'THEN
      IF (X=9) THEN 
        X<=0;
      ELSE 
        X<=X+1;
      END IF;
    END IF;
  END PROCESS;
  WITH X SELECT
    SAIDA_DISP<="1111110" WHEN 0,
                "0110000" WHEN 1,
                "1101101" WHEN 2,
                "1111001" WHEN 3,
                "0110011" WHEN 4,
                "1011011" WHEN 5,
                "1011111" WHEN 6,
                "1110000" WHEN 7,
                "1111111" WHEN 8,
                "1111011" WHEN 9;
END ONE;

ENTITY MUX IS
  PORT(
        CLK: IN BIT;
  DISPA,DISPV: IN BIT_VECTOR(6 DOWNTO 0);
  SAIDA_DISP: OUT BIT_VECTOR(6 DOWNTO 0);--A..G
  ENABLE_DISPA,ENABLE_DISPV:OUT BIT);
END MUX;

ARCHITECTURE ONE OF MUX IS
  SIGNAL X: INTEGER RANGE 0 TO 3:=0;
BEGIN
  PROCESS (CLK)
  BEGIN 
    IF  CLK'EVENT AND CLK='1'THEN
      IF (X=3) THEN 
        X<=0;
      ELSE 
        X<=X+1;
      END IF;
    END IF;
  END PROCESS;
  WITH X SELECT
    SAIDA_DISP<=DISPA WHEN 0,
                DISPV WHEN 1,
                DISPA WHEN 2,
                DISPV WHEN 3;

  WITH X SELECT
    ENABLE_DISPA<='1' WHEN 0,
                  '0' WHEN 1,
                  '1' WHEN 2,
                  '0'WHEN 3;
  WITH X SELECT
    ENABLE_DISPV<='0' WHEN 0,
                  '1' WHEN 1,
                  '0' WHEN 2,
                  '1' WHEN 3;			 
END ONE;
